//---------------------------------------------------------------------------
// Package: apb_pkg
//---------------------------------------------------------------------------
`ifndef APB_PKG
`define APB_PKG

`include "apb_define.sv"
`include "../ENV/apb_interface.sv"

package apb_pkg;
    import uvm_pkg::*;
    `include "uvm_macros.svh"

    `include "../ENV/apb_transaction.sv" 
    `include "../RAL/apb_reg_model.sv" 
    `include "../RAL/apb_reg_adapter.sv" 
    `include "../RAL/apb_reg_predictor.sv" 
    `include "../ENV/apb_sequence.sv" 
    `include "../ENV/apb_sequencer.sv" 
    `include "../ENV/apb_driver.sv" 
    `include "../ENV/apb_monitor.sv" 
    `include "../ENV/apb_agent.sv" 
    `include "../ENV/apb_env.sv" 
    `include "../TEST/apb_base_test.sv" 
    `include "../TEST/apb_sanity_test.sv" 
    `include "../TEST/apb_reg_test.sv" 
endpackage

`endif
