//---------------------------------------------------------------------------
// Defines: apb_define
//---------------------------------------------------------------------------
`define ADDRWIDTH 32
`define DATAWIDTH 32

`define IN_SKEW 0     // Clocking block skew to avoid setup violation
`define OUT_SKEW 0    // Clocking block skew to avoid hold violation
