//---------------------------------------------------------------------------
// uvm_reg_predictor Class: apb_reg_predictor
//---------------------------------------------------------------------------
`ifndef APB_REG_PREDICTOR
`define APB_REG_PREDICTOR

typedef uvm_reg_predictor#(apb_transaction) apb_reg_predictor;

`endif
